module main

import tf

fn main() {
	println(tf.version())
}