module main

import tf

fn main() {
	graph := tf.new_graph()

	graph.delete()
}