module main

import tf 

fn main() {
	s := tf.string_from("Hello Tf from V")

	println("stringify(s) = ${s.str()}")
}