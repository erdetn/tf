module main

import tf

fn main() {
	tf_code := tf.Code(6)

	println(tf_code.str())
}
